`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        //  $readmemh("code.mem", rom);
    //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _ op // R-Type
    // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1
    // rom[1] = 32'b0100000_00001_00010_000_00101_0110011;// sub x5, x2, x1
    // rom[2] = 32'b0000000_00000_00011_111_00110_0110011;// and x6, x3, x0
    // rom[3] = 32'b0000000_00000_00011_110_00111_0110011;// or  x7, x3, x0
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // rom[4] = 32'b0000000_00010_00000_010_01000_0100011;// sw x2, 8(x0)
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // B-Type
    // rom[5] = 32'b0000000_00010_00010_000_01100_1100011;// beq x2, x2, 12
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    // rom[6] = 32'b000000001000_00000_010_01000_0000011;// lw x8, 8(x0)
    
    
    // rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
// //   ... existing code ...
//     rom[0] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1 
//     rom[1] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4 
//     rom[2] = 32'b000000000001_00010_110_01011_0010011;// ori x11, x2, 1 
//     rom[3] = 32'b000000000011_00001_001_01100_0010011;// slli x12, x1, 3
//     rom[4] = 32'b000000000010_00001_010_01101_0010011;// slti x13, x1, 2
//     rom[5] = 32'b000000000011_00001_011_01110_0010011;// sltiu x14, x1, 3
//     rom[6] = 32'b000000000101_00001_100_01111_0010011;// xori x15, x1, 5
//     rom[7] = 32'b000000000010_00001_101_10000_0010011;// srli x16, x1, 2
//     rom[8] = 32'b010000000010_00001_101_10001_0010011;// srai x17, x1, 2
// //... existing code ...

//... existing code ...
    // Load/Store 부호 확장 테스트 시퀀스
    rom[0] = 32'b111111111111_00001_000_01001_0010011;// addi x9, x1, -1    // x9 = 0 (1-1)
    rom[1] = 32'b111111111110_00001_000_01010_0010011;// addi x10, x1, -2   // x10 = -1 (1-2)
    rom[2] = 32'b111111111101_00001_000_01011_0010011;// addi x11, x1, -3   // x11 = -2 (1-3)
    rom[3] = 32'b111111111100_00001_000_01100_0010011;// addi x12, x1, -4   // x12 = -3 (1-4)
    
    // Store 명령어들 - 음수 값들을 저장
    rom[4] = 32'b0000000_01010_00000_000_00100_0100011;// sb x10, 4(x0)     // Store byte -1 at addr 4
    rom[5] = 32'b0000000_01011_00000_001_00110_0100011;// sh x11, 6(x0)     // Store halfword -2 at addr 6
    rom[6] = 32'b0000000_01100_00000_010_01000_0100011;// sw x12, 8(x0)     // Store word -3 at addr 8
    
    // Load 명령어들 - 부호 확장 차이 확인
    rom[7] = 32'b000000000100_00000_000_01101_0000011;// lb x13, 4(x0)      // Load signed byte: -1 (부호 확장)
    rom[8] = 32'b000000000110_00000_001_01110_0000011;// lh x14, 6(x0)      // Load signed halfword: -2 (부호 확장)
    rom[9] = 32'b000000001000_00000_010_01111_0000011;// lw x15, 8(x0)      // Load word: -3
    rom[10] = 32'b000000000100_00000_100_10000_0000011;// lbu x16, 4(x0)     // Load unsigned byte: 255 (부호 확장 없음)
    rom[11] = 32'b000000000110_00000_101_10001_0000011;// lhu x17, 6(x0)     // Load unsigned halfword: 65534 (부호 확장 없음)
// ... existing code ...

  
    // second check
    // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1
    // rom[1] = 32'b0100000_00001_00010_000_00101_0110011;// sub x5, x2, x1
    // rom[2] = 32'b0000000_00000_00011_111_00110_0110011;// and x6, x3, x0
    // rom[3] = 32'b0000000_00000_00011_110_00111_0110011;// or  x7, x3, x0
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // S-Type
    // rom[0] = 32'b0000000_00001_00000_010_01000_0100011;// sw x1, 8(x0)
    // rom[1] = 32'b0000000_00010_00000_000_01011_0100011;// sb x2, 11(x0) - Store Byte
    //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ op // B-Type
    // rom[6] = 32'b0000000_00010_00010_000_01100_1100011;// beq x2, x2, 12
    //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // L-Type
    // rom[0] = 32'b000000000000_00000_010_00001_0000011;// lw x1, 8(x0)
    // rom[0] = 32'b0000000_00001_00000_000_00001_0100011;// sb x1, 1(x0)
    // rom[1] = 32'b000000000001_00000_000_00001_0000011;// lb x1, 1(x0)
    // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ op // I-Type
    // rom[8] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1 
    // rom[9] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4 
    // rom[10] = 32'b000000000001_00010_110_01011_0010011;// ori x11, x2, 1 
    // rom[11] = 32'b000000000011_00001_001_01100_0010011;// slli x12, x1, 1 // 2b00001011 << 3 
    end

    assign data = rom[addr[31:2]];
endmodule
